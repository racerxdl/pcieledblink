// pcie2ram.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module pcie2ram (
		input  wire        clk_clk,                 //            clk.clk
		output wire        clk_125_clk,             //        clk_125.clk
		input  wire [31:0] hip_ctrl_test_in,        //       hip_ctrl.test_in
		input  wire        hip_ctrl_simu_mode_pipe, //               .simu_mode_pipe
		input  wire        hip_npor_npor,           //       hip_npor.npor
		input  wire        hip_npor_pin_perst,      //               .pin_perst
		input  wire        hip_refclk_clk,          //     hip_refclk.clk
		input  wire        hip_serial_rx_in0,       //     hip_serial.rx_in0
		output wire        hip_serial_tx_out0,      //               .tx_out0
		input  wire [11:0] pcie_ram_bus_address,    //   pcie_ram_bus.address
		input  wire        pcie_ram_bus_chipselect, //               .chipselect
		input  wire        pcie_ram_bus_clken,      //               .clken
		input  wire        pcie_ram_bus_write,      //               .write
		output wire [63:0] pcie_ram_bus_readdata,   //               .readdata
		input  wire [63:0] pcie_ram_bus_writedata,  //               .writedata
		input  wire [7:0]  pcie_ram_bus_byteenable, //               .byteenable
		input  wire        pcie_ram_clk_clk,        //   pcie_ram_clk.clk
		input  wire        pcie_ram_reset_reset,    // pcie_ram_reset.reset
		input  wire        reset_reset_n            //          reset.reset_n
	);

	wire          pcie_hip_coreclkout_clk;                               // pcie_hip:coreclkout -> [mm_interconnect_0:pcie_hip_coreclkout_clk, pcie_ram:clk, rst_controller:clk]
	wire   [91:0] pcie_hip_reconfig_from_xcvr_reconfig_from_xcvr;        // pcie_hip:reconfig_from_xcvr -> pcie_reconfig:reconfig_from_xcvr
	wire  [139:0] pcie_reconfig_reconfig_to_xcvr_reconfig_to_xcvr;       // pcie_reconfig:reconfig_to_xcvr -> pcie_hip:reconfig_to_xcvr
	wire          pcie_hip_rxm_bar0_waitrequest;                         // mm_interconnect_0:pcie_hip_Rxm_BAR0_waitrequest -> pcie_hip:RxmWaitRequest_0_i
	wire   [63:0] pcie_hip_rxm_bar0_readdata;                            // mm_interconnect_0:pcie_hip_Rxm_BAR0_readdata -> pcie_hip:RxmReadData_0_i
	wire   [31:0] pcie_hip_rxm_bar0_address;                             // pcie_hip:RxmAddress_0_o -> mm_interconnect_0:pcie_hip_Rxm_BAR0_address
	wire          pcie_hip_rxm_bar0_read;                                // pcie_hip:RxmRead_0_o -> mm_interconnect_0:pcie_hip_Rxm_BAR0_read
	wire    [7:0] pcie_hip_rxm_bar0_byteenable;                          // pcie_hip:RxmByteEnable_0_o -> mm_interconnect_0:pcie_hip_Rxm_BAR0_byteenable
	wire          pcie_hip_rxm_bar0_readdatavalid;                       // mm_interconnect_0:pcie_hip_Rxm_BAR0_readdatavalid -> pcie_hip:RxmReadDataValid_0_i
	wire          pcie_hip_rxm_bar0_write;                               // pcie_hip:RxmWrite_0_o -> mm_interconnect_0:pcie_hip_Rxm_BAR0_write
	wire   [63:0] pcie_hip_rxm_bar0_writedata;                           // pcie_hip:RxmWriteData_0_o -> mm_interconnect_0:pcie_hip_Rxm_BAR0_writedata
	wire    [6:0] pcie_hip_rxm_bar0_burstcount;                          // pcie_hip:RxmBurstCount_0_o -> mm_interconnect_0:pcie_hip_Rxm_BAR0_burstcount
	wire   [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata; // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire    [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;  // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire          mm_interconnect_0_pcie_ram_s1_chipselect;              // mm_interconnect_0:pcie_ram_s1_chipselect -> pcie_ram:chipselect
	wire  [127:0] mm_interconnect_0_pcie_ram_s1_readdata;                // pcie_ram:readdata -> mm_interconnect_0:pcie_ram_s1_readdata
	wire   [10:0] mm_interconnect_0_pcie_ram_s1_address;                 // mm_interconnect_0:pcie_ram_s1_address -> pcie_ram:address
	wire   [15:0] mm_interconnect_0_pcie_ram_s1_byteenable;              // mm_interconnect_0:pcie_ram_s1_byteenable -> pcie_ram:byteenable
	wire          mm_interconnect_0_pcie_ram_s1_write;                   // mm_interconnect_0:pcie_ram_s1_write -> pcie_ram:write
	wire  [127:0] mm_interconnect_0_pcie_ram_s1_writedata;               // mm_interconnect_0:pcie_ram_s1_writedata -> pcie_ram:writedata
	wire          mm_interconnect_0_pcie_ram_s1_clken;                   // mm_interconnect_0:pcie_ram_s1_clken -> pcie_ram:clken
	wire          rst_controller_reset_out_reset;                        // rst_controller:reset_out -> [mm_interconnect_0:pcie_ram_reset1_reset_bridge_in_reset_reset, pcie_ram:reset]
	wire          pcie_hip_nreset_status_reset;                          // pcie_hip:reset_status -> [rst_controller:reset_in0, rst_controller_002:reset_in0]
	wire          rst_controller_001_reset_out_reset;                    // rst_controller_001:reset_out -> pcie_reconfig:mgmt_rst_reset
	wire          rst_controller_002_reset_out_reset;                    // rst_controller_002:reset_out -> [mm_interconnect_0:sysid_qsys_0_reset_reset_bridge_in_reset_reset, sysid_qsys_0:reset_n]

	altpcie_sv_hip_avmm_hwtcl #(
		.lane_mask_hwtcl                          ("x1"),
		.gen123_lane_rate_mode_hwtcl              ("Gen1 (2.5 Gbps)"),
		.port_type_hwtcl                          ("Native endpoint"),
		.pcie_spec_version_hwtcl                  ("2.1"),
		.pll_refclk_freq_hwtcl                    ("100 MHz"),
		.set_pld_clk_x1_625MHz_hwtcl              (0),
		.in_cvp_mode_hwtcl                        (0),
		.enable_tl_only_sim_hwtcl                 (0),
		.use_atx_pll_hwtcl                        (0),
		.enable_power_on_rst_pulse_hwtcl          (0),
		.enable_pcisigtest_hwtcl                  (0),
		.bar0_size_mask_hwtcl                     (21),
		.bar0_io_space_hwtcl                      ("Disabled"),
		.bar0_64bit_mem_space_hwtcl               ("Disabled"),
		.bar0_prefetchable_hwtcl                  ("Disabled"),
		.bar1_size_mask_hwtcl                     (0),
		.bar1_io_space_hwtcl                      ("Disabled"),
		.bar1_prefetchable_hwtcl                  ("Disabled"),
		.bar2_size_mask_hwtcl                     (0),
		.bar2_io_space_hwtcl                      ("Disabled"),
		.bar2_64bit_mem_space_hwtcl               ("Disabled"),
		.bar2_prefetchable_hwtcl                  ("Disabled"),
		.bar3_size_mask_hwtcl                     (0),
		.bar3_io_space_hwtcl                      ("Disabled"),
		.bar3_prefetchable_hwtcl                  ("Disabled"),
		.bar4_size_mask_hwtcl                     (0),
		.bar4_io_space_hwtcl                      ("Disabled"),
		.bar4_64bit_mem_space_hwtcl               ("Disabled"),
		.bar4_prefetchable_hwtcl                  ("Disabled"),
		.bar5_size_mask_hwtcl                     (0),
		.bar5_io_space_hwtcl                      ("Disabled"),
		.bar5_prefetchable_hwtcl                  ("Disabled"),
		.vendor_id_hwtcl                          (4466),
		.device_id_hwtcl                          (167),
		.revision_id_hwtcl                        (1),
		.class_code_hwtcl                         (0),
		.subsystem_vendor_id_hwtcl                (418),
		.subsystem_device_id_hwtcl                (1),
		.max_payload_size_hwtcl                   (128),
		.extend_tag_field_hwtcl                   ("32"),
		.completion_timeout_hwtcl                 ("ABCD"),
		.enable_completion_timeout_disable_hwtcl  (1),
		.use_aer_hwtcl                            (1),
		.ecrc_check_capable_hwtcl                 (0),
		.ecrc_gen_capable_hwtcl                   (0),
		.use_crc_forwarding_hwtcl                 (0),
		.port_link_number_hwtcl                   (1),
		.dll_active_report_support_hwtcl          (0),
		.surprise_down_error_support_hwtcl        (0),
		.slotclkcfg_hwtcl                         (1),
		.msi_multi_message_capable_hwtcl          ("4"),
		.msi_64bit_addressing_capable_hwtcl       ("true"),
		.msi_masking_capable_hwtcl                ("false"),
		.msi_support_hwtcl                        ("true"),
		.enable_function_msix_support_hwtcl       (0),
		.msix_table_size_hwtcl                    (0),
		.msix_table_offset_hwtcl                  ("0"),
		.msix_table_bir_hwtcl                     (0),
		.msix_pba_offset_hwtcl                    ("0"),
		.msix_pba_bir_hwtcl                       (0),
		.enable_slot_register_hwtcl               (0),
		.slot_power_scale_hwtcl                   (0),
		.slot_power_limit_hwtcl                   (0),
		.slot_number_hwtcl                        (0),
		.endpoint_l0_latency_hwtcl                (0),
		.endpoint_l1_latency_hwtcl                (0),
		.vsec_id_hwtcl                            (4466),
		.vsec_rev_hwtcl                           (0),
		.user_id_hwtcl                            (0),
		.avmm_width_hwtcl                         (64),
		.AVALON_ADDR_WIDTH                        (32),
		.avmm_burst_width_hwtcl                   (7),
		.CB_PCIE_MODE                             (1),
		.CB_PCIE_RX_LITE                          (0),
		.CB_RXM_DATA_WIDTH                        (64),
		.CG_AVALON_S_ADDR_WIDTH                   (21),
		.CG_IMPL_CRA_AV_SLAVE_PORT                (0),
		.CG_ENABLE_ADVANCED_INTERRUPT             (0),
		.CG_ENABLE_A2P_INTERRUPT                  (0),
		.CB_A2P_ADDR_MAP_IS_FIXED                 (0),
		.CB_A2P_ADDR_MAP_NUM_ENTRIES              (2),
		.BYPASSS_A2P_TRANSLATION                  (0),
		.a2p_pass_thru_bits                       (20),
		.ast_width_hwtcl                          ("Avalon-ST 64-bit"),
		.use_ast_parity                           (0),
		.millisecond_cycle_count_hwtcl            (124250),
		.port_width_be_hwtcl                      (8),
		.port_width_data_hwtcl                    (64),
		.hip_reconfig_hwtcl                       (0),
		.expansion_base_address_register_hwtcl    (0),
		.prefetchable_mem_window_addr_width_hwtcl (0),
		.bypass_cdc_hwtcl                         ("false"),
		.enable_rx_buffer_checking_hwtcl          ("false"),
		.disable_link_x2_support_hwtcl            ("false"),
		.wrong_device_id_hwtcl                    ("disable"),
		.data_pack_rx_hwtcl                       ("disable"),
		.ltssm_1ms_timeout_hwtcl                  ("disable"),
		.ltssm_freqlocked_check_hwtcl             ("disable"),
		.deskew_comma_hwtcl                       ("skp_eieos_deskw"),
		.device_number_hwtcl                      (0),
		.pipex1_debug_sel_hwtcl                   ("disable"),
		.pclk_out_sel_hwtcl                       ("pclk"),
		.no_soft_reset_hwtcl                      ("false"),
		.maximum_current_hwtcl                    (0),
		.d1_support_hwtcl                         ("false"),
		.d2_support_hwtcl                         ("false"),
		.d0_pme_hwtcl                             ("false"),
		.d1_pme_hwtcl                             ("false"),
		.d2_pme_hwtcl                             ("false"),
		.d3_hot_pme_hwtcl                         ("false"),
		.d3_cold_pme_hwtcl                        ("false"),
		.low_priority_vc_hwtcl                    ("single_vc"),
		.disable_snoop_packet_hwtcl               ("false"),
		.enable_l1_aspm_hwtcl                     ("false"),
		.rx_ei_l0s_hwtcl                          (0),
		.enable_l0s_aspm_hwtcl                    ("false"),
		.aspm_config_management_hwtcl             ("true"),
		.l1_exit_latency_sameclock_hwtcl          (0),
		.l1_exit_latency_diffclock_hwtcl          (0),
		.hot_plug_support_hwtcl                   (0),
		.extended_tag_reset_hwtcl                 ("false"),
		.no_command_completed_hwtcl               ("false"),
		.interrupt_pin_hwtcl                      ("inta"),
		.bridge_port_vga_enable_hwtcl             ("false"),
		.bridge_port_ssid_support_hwtcl           ("false"),
		.ssvid_hwtcl                              (0),
		.ssid_hwtcl                               (0),
		.eie_before_nfts_count_hwtcl              (4),
		.gen2_diffclock_nfts_count_hwtcl          (255),
		.gen2_sameclock_nfts_count_hwtcl          (255),
		.l0_exit_latency_sameclock_hwtcl          (6),
		.l0_exit_latency_diffclock_hwtcl          (6),
		.atomic_op_routing_hwtcl                  ("false"),
		.atomic_op_completer_32bit_hwtcl          ("false"),
		.atomic_op_completer_64bit_hwtcl          ("false"),
		.cas_completer_128bit_hwtcl               ("false"),
		.ltr_mechanism_hwtcl                      ("false"),
		.tph_completer_hwtcl                      ("false"),
		.extended_format_field_hwtcl              ("false"),
		.atomic_malformed_hwtcl                   ("true"),
		.flr_capability_hwtcl                     ("false"),
		.enable_adapter_half_rate_mode_hwtcl      ("false"),
		.vc0_clk_enable_hwtcl                     ("true"),
		.register_pipe_signals_hwtcl              ("false"),
		.skp_os_gen3_count_hwtcl                  (0),
		.tx_cdc_almost_empty_hwtcl                (5),
		.rx_l0s_count_idl_hwtcl                   (0),
		.cdc_dummy_insert_limit_hwtcl             (11),
		.ei_delay_powerdown_count_hwtcl           (10),
		.skp_os_schedule_count_hwtcl              (0),
		.fc_init_timer_hwtcl                      (1024),
		.l01_entry_latency_hwtcl                  (31),
		.flow_control_update_count_hwtcl          (30),
		.flow_control_timeout_count_hwtcl         (200),
		.retry_buffer_last_active_address_hwtcl   (2047),
		.reserved_debug_hwtcl                     (0),
		.bypass_clk_switch_hwtcl                  ("false"),
		.l2_async_logic_hwtcl                     ("disable"),
		.indicator_hwtcl                          (0),
		.diffclock_nfts_count_hwtcl               (128),
		.sameclock_nfts_count_hwtcl               (128),
		.rx_cdc_almost_full_hwtcl                 (12),
		.tx_cdc_almost_full_hwtcl                 (11),
		.credit_buffer_allocation_aux_hwtcl       ("absolute"),
		.vc0_rx_flow_ctrl_posted_header_hwtcl     (16),
		.vc0_rx_flow_ctrl_posted_data_hwtcl       (16),
		.vc0_rx_flow_ctrl_nonposted_header_hwtcl  (16),
		.vc0_rx_flow_ctrl_nonposted_data_hwtcl    (0),
		.vc0_rx_flow_ctrl_compl_header_hwtcl      (0),
		.vc0_rx_flow_ctrl_compl_data_hwtcl        (0),
		.cpl_spc_header_hwtcl                     (195),
		.cpl_spc_data_hwtcl                       (781),
		.gen3_rxfreqlock_counter_hwtcl            (0),
		.gen3_skip_ph2_ph3_hwtcl                  (0),
		.g3_bypass_equlz_hwtcl                    (0),
		.cvp_data_compressed_hwtcl                ("false"),
		.cvp_data_encrypted_hwtcl                 ("false"),
		.cvp_mode_reset_hwtcl                     ("false"),
		.cvp_clk_reset_hwtcl                      ("false"),
		.cseb_cpl_status_during_cvp_hwtcl         ("completer_abort"),
		.core_clk_sel_hwtcl                       ("core_clk_250"),
		.cvp_rate_sel_hwtcl                       ("full_rate"),
		.g3_dis_rx_use_prst_hwtcl                 ("true"),
		.g3_dis_rx_use_prst_ep_hwtcl              ("true"),
		.deemphasis_enable_hwtcl                  ("false"),
		.reconfig_to_xcvr_width                   (140),
		.reconfig_from_xcvr_width                 (92),
		.single_rx_detect_hwtcl                   (1),
		.hip_hard_reset_hwtcl                     (1),
		.use_cvp_update_core_pof_hwtcl            (0),
		.pcie_inspector_hwtcl                     (0),
		.tlp_inspector_hwtcl                      (0),
		.tlp_inspector_use_signal_probe_hwtcl     (0),
		.tlp_insp_trg_dw0_hwtcl                   (2049),
		.tlp_insp_trg_dw1_hwtcl                   (0),
		.tlp_insp_trg_dw2_hwtcl                   (0),
		.tlp_insp_trg_dw3_hwtcl                   (0),
		.hwtcl_override_g2_txvod                  (1),
		.rpre_emph_a_val_hwtcl                    (9),
		.rpre_emph_b_val_hwtcl                    (0),
		.rpre_emph_c_val_hwtcl                    (16),
		.rpre_emph_d_val_hwtcl                    (13),
		.rpre_emph_e_val_hwtcl                    (5),
		.rvod_sel_a_val_hwtcl                     (42),
		.rvod_sel_b_val_hwtcl                     (38),
		.rvod_sel_c_val_hwtcl                     (38),
		.rvod_sel_d_val_hwtcl                     (43),
		.rvod_sel_e_val_hwtcl                     (15)
	) pcie_hip (
		.coreclkout           (pcie_hip_coreclkout_clk),                         //          coreclkout.clk
		.refclk               (hip_refclk_clk),                                  //              refclk.clk
		.npor                 (hip_npor_npor),                                   //                npor.npor
		.pin_perst            (hip_npor_pin_perst),                              //                    .pin_perst
		.reset_status         (pcie_hip_nreset_status_reset),                    //       nreset_status.reset_n
		.RxmAddress_0_o       (pcie_hip_rxm_bar0_address),                       //            Rxm_BAR0.address
		.RxmRead_0_o          (pcie_hip_rxm_bar0_read),                          //                    .read
		.RxmWaitRequest_0_i   (pcie_hip_rxm_bar0_waitrequest),                   //                    .waitrequest
		.RxmWrite_0_o         (pcie_hip_rxm_bar0_write),                         //                    .write
		.RxmReadDataValid_0_i (pcie_hip_rxm_bar0_readdatavalid),                 //                    .readdatavalid
		.RxmReadData_0_i      (pcie_hip_rxm_bar0_readdata),                      //                    .readdata
		.RxmWriteData_0_o     (pcie_hip_rxm_bar0_writedata),                     //                    .writedata
		.RxmBurstCount_0_o    (pcie_hip_rxm_bar0_burstcount),                    //                    .burstcount
		.RxmByteEnable_0_o    (pcie_hip_rxm_bar0_byteenable),                    //                    .byteenable
		.derr_cor_ext_rcv     (),                                                //          hip_status.derr_cor_ext_rcv
		.derr_cor_ext_rpl     (),                                                //                    .derr_cor_ext_rpl
		.derr_rpl             (),                                                //                    .derr_rpl
		.dlup                 (),                                                //                    .dlup
		.dlup_exit            (),                                                //                    .dlup_exit
		.ev128ns              (),                                                //                    .ev128ns
		.ev1us                (),                                                //                    .ev1us
		.hotrst_exit          (),                                                //                    .hotrst_exit
		.int_status           (),                                                //                    .int_status
		.l2_exit              (),                                                //                    .l2_exit
		.lane_act             (),                                                //                    .lane_act
		.ltssmstate           (),                                                //                    .ltssmstate
		.rx_par_err           (),                                                //                    .rx_par_err
		.tx_par_err           (),                                                //                    .tx_par_err
		.cfg_par_err          (),                                                //                    .cfg_par_err
		.ko_cpl_spc_header    (),                                                //                    .ko_cpl_spc_header
		.ko_cpl_spc_data      (),                                                //                    .ko_cpl_spc_data
		.currentspeed         (),                                                //    hip_currentspeed.currentspeed
		.reconfig_to_xcvr     (pcie_reconfig_reconfig_to_xcvr_reconfig_to_xcvr), //    reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr   (pcie_hip_reconfig_from_xcvr_reconfig_from_xcvr),  //  reconfig_from_xcvr.reconfig_from_xcvr
		.fixedclk_locked      (),                                                // reconfig_clk_locked.fixedclk_locked
		.rx_in0               (hip_serial_rx_in0),                               //          hip_serial.rx_in0
		.tx_out0              (hip_serial_tx_out0),                              //                    .tx_out0
		.sim_pipe_pclk_in     (),                                                //            hip_pipe.sim_pipe_pclk_in
		.sim_pipe_rate        (),                                                //                    .sim_pipe_rate
		.sim_ltssmstate       (),                                                //                    .sim_ltssmstate
		.eidleinfersel0       (),                                                //                    .eidleinfersel0
		.powerdown0           (),                                                //                    .powerdown0
		.rxpolarity0          (),                                                //                    .rxpolarity0
		.txcompl0             (),                                                //                    .txcompl0
		.txdata0              (),                                                //                    .txdata0
		.txdatak0             (),                                                //                    .txdatak0
		.txdetectrx0          (),                                                //                    .txdetectrx0
		.txelecidle0          (),                                                //                    .txelecidle0
		.txdeemph0            (),                                                //                    .txdeemph0
		.txmargin0            (),                                                //                    .txmargin0
		.txswing0             (),                                                //                    .txswing0
		.phystatus0           (),                                                //                    .phystatus0
		.rxdata0              (),                                                //                    .rxdata0
		.rxdatak0             (),                                                //                    .rxdatak0
		.rxelecidle0          (),                                                //                    .rxelecidle0
		.rxstatus0            (),                                                //                    .rxstatus0
		.rxvalid0             (),                                                //                    .rxvalid0
		.test_in              (hip_ctrl_test_in),                                //            hip_ctrl.test_in
		.simu_mode_pipe       (hip_ctrl_simu_mode_pipe),                         //                    .simu_mode_pipe
		.rx_in1               (1'b0),                                            //         (terminated)
		.rx_in2               (1'b0),                                            //         (terminated)
		.rx_in3               (1'b0),                                            //         (terminated)
		.rx_in4               (1'b0),                                            //         (terminated)
		.rx_in5               (1'b0),                                            //         (terminated)
		.rx_in6               (1'b0),                                            //         (terminated)
		.rx_in7               (1'b0),                                            //         (terminated)
		.tx_out1              (),                                                //         (terminated)
		.tx_out2              (),                                                //         (terminated)
		.tx_out3              (),                                                //         (terminated)
		.tx_out4              (),                                                //         (terminated)
		.tx_out5              (),                                                //         (terminated)
		.tx_out6              (),                                                //         (terminated)
		.tx_out7              (),                                                //         (terminated)
		.eidleinfersel1       (),                                                //         (terminated)
		.eidleinfersel2       (),                                                //         (terminated)
		.eidleinfersel3       (),                                                //         (terminated)
		.eidleinfersel4       (),                                                //         (terminated)
		.eidleinfersel5       (),                                                //         (terminated)
		.eidleinfersel6       (),                                                //         (terminated)
		.eidleinfersel7       (),                                                //         (terminated)
		.powerdown1           (),                                                //         (terminated)
		.powerdown2           (),                                                //         (terminated)
		.powerdown3           (),                                                //         (terminated)
		.powerdown4           (),                                                //         (terminated)
		.powerdown5           (),                                                //         (terminated)
		.powerdown6           (),                                                //         (terminated)
		.powerdown7           (),                                                //         (terminated)
		.rxpolarity1          (),                                                //         (terminated)
		.rxpolarity2          (),                                                //         (terminated)
		.rxpolarity3          (),                                                //         (terminated)
		.rxpolarity4          (),                                                //         (terminated)
		.rxpolarity5          (),                                                //         (terminated)
		.rxpolarity6          (),                                                //         (terminated)
		.rxpolarity7          (),                                                //         (terminated)
		.txcompl1             (),                                                //         (terminated)
		.txcompl2             (),                                                //         (terminated)
		.txcompl3             (),                                                //         (terminated)
		.txcompl4             (),                                                //         (terminated)
		.txcompl5             (),                                                //         (terminated)
		.txcompl6             (),                                                //         (terminated)
		.txcompl7             (),                                                //         (terminated)
		.txdata1              (),                                                //         (terminated)
		.txdata2              (),                                                //         (terminated)
		.txdata3              (),                                                //         (terminated)
		.txdata4              (),                                                //         (terminated)
		.txdata5              (),                                                //         (terminated)
		.txdata6              (),                                                //         (terminated)
		.txdata7              (),                                                //         (terminated)
		.txdatak1             (),                                                //         (terminated)
		.txdatak2             (),                                                //         (terminated)
		.txdatak3             (),                                                //         (terminated)
		.txdatak4             (),                                                //         (terminated)
		.txdatak5             (),                                                //         (terminated)
		.txdatak6             (),                                                //         (terminated)
		.txdatak7             (),                                                //         (terminated)
		.txdetectrx1          (),                                                //         (terminated)
		.txdetectrx2          (),                                                //         (terminated)
		.txdetectrx3          (),                                                //         (terminated)
		.txdetectrx4          (),                                                //         (terminated)
		.txdetectrx5          (),                                                //         (terminated)
		.txdetectrx6          (),                                                //         (terminated)
		.txdetectrx7          (),                                                //         (terminated)
		.txelecidle1          (),                                                //         (terminated)
		.txelecidle2          (),                                                //         (terminated)
		.txelecidle3          (),                                                //         (terminated)
		.txelecidle4          (),                                                //         (terminated)
		.txelecidle5          (),                                                //         (terminated)
		.txelecidle6          (),                                                //         (terminated)
		.txelecidle7          (),                                                //         (terminated)
		.txdeemph1            (),                                                //         (terminated)
		.txdeemph2            (),                                                //         (terminated)
		.txdeemph3            (),                                                //         (terminated)
		.txdeemph4            (),                                                //         (terminated)
		.txdeemph5            (),                                                //         (terminated)
		.txdeemph6            (),                                                //         (terminated)
		.txdeemph7            (),                                                //         (terminated)
		.txmargin1            (),                                                //         (terminated)
		.txmargin2            (),                                                //         (terminated)
		.txmargin3            (),                                                //         (terminated)
		.txmargin4            (),                                                //         (terminated)
		.txmargin5            (),                                                //         (terminated)
		.txmargin6            (),                                                //         (terminated)
		.txmargin7            (),                                                //         (terminated)
		.txswing1             (),                                                //         (terminated)
		.txswing2             (),                                                //         (terminated)
		.txswing3             (),                                                //         (terminated)
		.txswing4             (),                                                //         (terminated)
		.txswing5             (),                                                //         (terminated)
		.txswing6             (),                                                //         (terminated)
		.txswing7             (),                                                //         (terminated)
		.phystatus1           (1'b0),                                            //         (terminated)
		.phystatus2           (1'b0),                                            //         (terminated)
		.phystatus3           (1'b0),                                            //         (terminated)
		.phystatus4           (1'b0),                                            //         (terminated)
		.phystatus5           (1'b0),                                            //         (terminated)
		.phystatus6           (1'b0),                                            //         (terminated)
		.phystatus7           (1'b0),                                            //         (terminated)
		.rxdata1              (8'b00000000),                                     //         (terminated)
		.rxdata2              (8'b00000000),                                     //         (terminated)
		.rxdata3              (8'b00000000),                                     //         (terminated)
		.rxdata4              (8'b00000000),                                     //         (terminated)
		.rxdata5              (8'b00000000),                                     //         (terminated)
		.rxdata6              (8'b00000000),                                     //         (terminated)
		.rxdata7              (8'b00000000),                                     //         (terminated)
		.rxdatak1             (1'b0),                                            //         (terminated)
		.rxdatak2             (1'b0),                                            //         (terminated)
		.rxdatak3             (1'b0),                                            //         (terminated)
		.rxdatak4             (1'b0),                                            //         (terminated)
		.rxdatak5             (1'b0),                                            //         (terminated)
		.rxdatak6             (1'b0),                                            //         (terminated)
		.rxdatak7             (1'b0),                                            //         (terminated)
		.rxelecidle1          (1'b0),                                            //         (terminated)
		.rxelecidle2          (1'b0),                                            //         (terminated)
		.rxelecidle3          (1'b0),                                            //         (terminated)
		.rxelecidle4          (1'b0),                                            //         (terminated)
		.rxelecidle5          (1'b0),                                            //         (terminated)
		.rxelecidle6          (1'b0),                                            //         (terminated)
		.rxelecidle7          (1'b0),                                            //         (terminated)
		.rxstatus1            (3'b000),                                          //         (terminated)
		.rxstatus2            (3'b000),                                          //         (terminated)
		.rxstatus3            (3'b000),                                          //         (terminated)
		.rxstatus4            (3'b000),                                          //         (terminated)
		.rxstatus5            (3'b000),                                          //         (terminated)
		.rxstatus6            (3'b000),                                          //         (terminated)
		.rxstatus7            (3'b000),                                          //         (terminated)
		.rxvalid1             (1'b0),                                            //         (terminated)
		.rxvalid2             (1'b0),                                            //         (terminated)
		.rxvalid3             (1'b0),                                            //         (terminated)
		.rxvalid4             (1'b0),                                            //         (terminated)
		.rxvalid5             (1'b0),                                            //         (terminated)
		.rxvalid6             (1'b0),                                            //         (terminated)
		.rxvalid7             (1'b0),                                            //         (terminated)
		.rxdataskip0          (1'b0),                                            //         (terminated)
		.rxdataskip1          (1'b0),                                            //         (terminated)
		.rxdataskip2          (1'b0),                                            //         (terminated)
		.rxdataskip3          (1'b0),                                            //         (terminated)
		.rxdataskip4          (1'b0),                                            //         (terminated)
		.rxdataskip5          (1'b0),                                            //         (terminated)
		.rxdataskip6          (1'b0),                                            //         (terminated)
		.rxdataskip7          (1'b0),                                            //         (terminated)
		.rxblkst0             (1'b0),                                            //         (terminated)
		.rxblkst1             (1'b0),                                            //         (terminated)
		.rxblkst2             (1'b0),                                            //         (terminated)
		.rxblkst3             (1'b0),                                            //         (terminated)
		.rxblkst4             (1'b0),                                            //         (terminated)
		.rxblkst5             (1'b0),                                            //         (terminated)
		.rxblkst6             (1'b0),                                            //         (terminated)
		.rxblkst7             (1'b0),                                            //         (terminated)
		.rxsynchd0            (2'b00),                                           //         (terminated)
		.rxsynchd1            (2'b00),                                           //         (terminated)
		.rxsynchd2            (2'b00),                                           //         (terminated)
		.rxsynchd3            (2'b00),                                           //         (terminated)
		.rxsynchd4            (2'b00),                                           //         (terminated)
		.rxsynchd5            (2'b00),                                           //         (terminated)
		.rxsynchd6            (2'b00),                                           //         (terminated)
		.rxsynchd7            (2'b00),                                           //         (terminated)
		.rxfreqlocked0        (1'b0),                                            //         (terminated)
		.rxfreqlocked1        (1'b0),                                            //         (terminated)
		.rxfreqlocked2        (1'b0),                                            //         (terminated)
		.rxfreqlocked3        (1'b0),                                            //         (terminated)
		.rxfreqlocked4        (1'b0),                                            //         (terminated)
		.rxfreqlocked5        (1'b0),                                            //         (terminated)
		.rxfreqlocked6        (1'b0),                                            //         (terminated)
		.rxfreqlocked7        (1'b0),                                            //         (terminated)
		.currentcoeff0        (),                                                //         (terminated)
		.currentcoeff1        (),                                                //         (terminated)
		.currentcoeff2        (),                                                //         (terminated)
		.currentcoeff3        (),                                                //         (terminated)
		.currentcoeff4        (),                                                //         (terminated)
		.currentcoeff5        (),                                                //         (terminated)
		.currentcoeff6        (),                                                //         (terminated)
		.currentcoeff7        (),                                                //         (terminated)
		.currentrxpreset0     (),                                                //         (terminated)
		.currentrxpreset1     (),                                                //         (terminated)
		.currentrxpreset2     (),                                                //         (terminated)
		.currentrxpreset3     (),                                                //         (terminated)
		.currentrxpreset4     (),                                                //         (terminated)
		.currentrxpreset5     (),                                                //         (terminated)
		.currentrxpreset6     (),                                                //         (terminated)
		.currentrxpreset7     (),                                                //         (terminated)
		.txsynchd0            (),                                                //         (terminated)
		.txsynchd1            (),                                                //         (terminated)
		.txsynchd2            (),                                                //         (terminated)
		.txsynchd3            (),                                                //         (terminated)
		.txsynchd4            (),                                                //         (terminated)
		.txsynchd5            (),                                                //         (terminated)
		.txsynchd6            (),                                                //         (terminated)
		.txsynchd7            (),                                                //         (terminated)
		.txblkst0             (),                                                //         (terminated)
		.txblkst1             (),                                                //         (terminated)
		.txblkst2             (),                                                //         (terminated)
		.txblkst3             (),                                                //         (terminated)
		.txblkst4             (),                                                //         (terminated)
		.txblkst5             (),                                                //         (terminated)
		.txblkst6             (),                                                //         (terminated)
		.txblkst7             ()                                                 //         (terminated)
	);

	pcie2ram_pcie_ram pcie_ram (
		.clk         (pcie_hip_coreclkout_clk),                  //   clk1.clk
		.address     (mm_interconnect_0_pcie_ram_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_pcie_ram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_pcie_ram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_pcie_ram_s1_write),      //       .write
		.readdata    (mm_interconnect_0_pcie_ram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_pcie_ram_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_pcie_ram_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),           // reset1.reset
		.address2    (pcie_ram_bus_address),                     //     s2.address
		.chipselect2 (pcie_ram_bus_chipselect),                  //       .chipselect
		.clken2      (pcie_ram_bus_clken),                       //       .clken
		.write2      (pcie_ram_bus_write),                       //       .write
		.readdata2   (pcie_ram_bus_readdata),                    //       .readdata
		.writedata2  (pcie_ram_bus_writedata),                   //       .writedata
		.byteenable2 (pcie_ram_bus_byteenable),                  //       .byteenable
		.clk2        (pcie_ram_clk_clk),                         //   clk2.clk
		.reset2      (pcie_ram_reset_reset),                     // reset2.reset
		.reset_req   (1'b0),                                     // (terminated)
		.freeze      (1'b0),                                     // (terminated)
		.reset_req2  (1'b0)                                      // (terminated)
	);

	alt_xcvr_reconfig #(
		.device_family                 ("Stratix V"),
		.number_of_reconfig_interfaces (2),
		.enable_offset                 (1),
		.enable_lc                     (1),
		.enable_dcd                    (0),
		.enable_dcd_power_up           (1),
		.enable_analog                 (0),
		.enable_eyemon                 (0),
		.enable_ber                    (0),
		.enable_dfe                    (0),
		.enable_adce                   (0),
		.enable_mif                    (0),
		.enable_pll                    (0)
	) pcie_reconfig (
		.reconfig_busy             (),                                                //      reconfig_busy.reconfig_busy
		.mgmt_clk_clk              (clk_clk),                                         //       mgmt_clk_clk.clk
		.mgmt_rst_reset            (rst_controller_001_reset_out_reset),              //     mgmt_rst_reset.reset
		.reconfig_mgmt_address     (),                                                //      reconfig_mgmt.address
		.reconfig_mgmt_read        (),                                                //                   .read
		.reconfig_mgmt_readdata    (),                                                //                   .readdata
		.reconfig_mgmt_waitrequest (),                                                //                   .waitrequest
		.reconfig_mgmt_write       (),                                                //                   .write
		.reconfig_mgmt_writedata   (),                                                //                   .writedata
		.reconfig_to_xcvr          (pcie_reconfig_reconfig_to_xcvr_reconfig_to_xcvr), //   reconfig_to_xcvr.reconfig_to_xcvr
		.reconfig_from_xcvr        (pcie_hip_reconfig_from_xcvr_reconfig_from_xcvr),  // reconfig_from_xcvr.reconfig_from_xcvr
		.tx_cal_busy               (),                                                //        (terminated)
		.rx_cal_busy               (),                                                //        (terminated)
		.cal_busy_in               (1'b0),                                            //        (terminated)
		.reconfig_mif_address      (),                                                //        (terminated)
		.reconfig_mif_read         (),                                                //        (terminated)
		.reconfig_mif_readdata     (16'b0000000000000000),                            //        (terminated)
		.reconfig_mif_waitrequest  (1'b0)                                             //        (terminated)
	);

	pcie2ram_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	pcie2ram_mm_interconnect_0 mm_interconnect_0 (
		.clk_125_clk_clk                                (clk_clk),                                               //                              clk_125_clk.clk
		.pcie_hip_coreclkout_clk                        (pcie_hip_coreclkout_clk),                               //                      pcie_hip_coreclkout.clk
		.pcie_ram_reset1_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                        //    pcie_ram_reset1_reset_bridge_in_reset.reset
		.sysid_qsys_0_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                    // sysid_qsys_0_reset_reset_bridge_in_reset.reset
		.pcie_hip_Rxm_BAR0_address                      (pcie_hip_rxm_bar0_address),                             //                        pcie_hip_Rxm_BAR0.address
		.pcie_hip_Rxm_BAR0_waitrequest                  (pcie_hip_rxm_bar0_waitrequest),                         //                                         .waitrequest
		.pcie_hip_Rxm_BAR0_burstcount                   (pcie_hip_rxm_bar0_burstcount),                          //                                         .burstcount
		.pcie_hip_Rxm_BAR0_byteenable                   (pcie_hip_rxm_bar0_byteenable),                          //                                         .byteenable
		.pcie_hip_Rxm_BAR0_read                         (pcie_hip_rxm_bar0_read),                                //                                         .read
		.pcie_hip_Rxm_BAR0_readdata                     (pcie_hip_rxm_bar0_readdata),                            //                                         .readdata
		.pcie_hip_Rxm_BAR0_readdatavalid                (pcie_hip_rxm_bar0_readdatavalid),                       //                                         .readdatavalid
		.pcie_hip_Rxm_BAR0_write                        (pcie_hip_rxm_bar0_write),                               //                                         .write
		.pcie_hip_Rxm_BAR0_writedata                    (pcie_hip_rxm_bar0_writedata),                           //                                         .writedata
		.pcie_ram_s1_address                            (mm_interconnect_0_pcie_ram_s1_address),                 //                              pcie_ram_s1.address
		.pcie_ram_s1_write                              (mm_interconnect_0_pcie_ram_s1_write),                   //                                         .write
		.pcie_ram_s1_readdata                           (mm_interconnect_0_pcie_ram_s1_readdata),                //                                         .readdata
		.pcie_ram_s1_writedata                          (mm_interconnect_0_pcie_ram_s1_writedata),               //                                         .writedata
		.pcie_ram_s1_byteenable                         (mm_interconnect_0_pcie_ram_s1_byteenable),              //                                         .byteenable
		.pcie_ram_s1_chipselect                         (mm_interconnect_0_pcie_ram_s1_chipselect),              //                                         .chipselect
		.pcie_ram_s1_clken                              (mm_interconnect_0_pcie_ram_s1_clken),                   //                                         .clken
		.sysid_qsys_0_control_slave_address             (mm_interconnect_0_sysid_qsys_0_control_slave_address),  //               sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata            (mm_interconnect_0_sysid_qsys_0_control_slave_readdata)  //                                         .readdata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~pcie_hip_nreset_status_reset),  // reset_in0.reset
		.clk            (pcie_hip_coreclkout_clk),        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~pcie_hip_nreset_status_reset),      // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	assign clk_125_clk = clk_clk;

endmodule
